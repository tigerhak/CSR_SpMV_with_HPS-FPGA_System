`timescale 1ns / 1ps

module tb_fp_dot;

	reg	[127:0]in_a;
	reg	[127:0]in_b;
	reg	clk, n_rst;
	wire	[31:0]out_c;
	
	fp_dot uut (
		.in_a(in_a),
		.in_b(in_b),
		.clk(clk),
		.n_rst(n_rst),
		.out_c(out_c)
	);

	initial begin
		clk = 0;
		n_rst = 0; #2000;
		n_rst = 1;
		in_a = 128'b00111111100000000000000000000000_01000000000000000000000000000000_01000000010000000000000000000000_01000000100000000000000000000000; 
		// (1, 2, 3, 4)
		in_b = 128'b01000000100000000000000000000000_01000000010000000000000000000000_01000000000000000000000000000000_00111111100000000000000000000000;
		// (4, 3, 2, 1)
		#100;
		
		in_a = 128'b00000000000000000000000000000000_01000000000000000000000000000000_00000000000000000000000000000000_01000100111110100000000000000000; 
		// (0, 2, 0, 2000)
		in_b = 128'b01000100011110100000000000000000_01000000010000000000000000000000_01000000000000000000000000000000_01000001001000000000000000000000;
		// (1000, 3, 2, 10)
		#100;
	end
     
	always #10 clk = !clk;
endmodule
